module IMEM (	
    input [29:0] PC_Out,
    output [31:0] instruction
);
    reg [31:0] memory [0:1023];
    assign instruction = memory[addr];
endmodule 
